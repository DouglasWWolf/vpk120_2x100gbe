//====================================================================================
//                        ------->  Revision History  <------
//====================================================================================
//
//   Date     Who   Ver  Changes
//====================================================================================
// 15-Aug-24  DWW     1  Initial creation
//====================================================================================

/*
     This module provides configuration for the downstream "packet generator"
*/


module packet_config # (parameter AW=8, parameter DEFAULT_INIT_VALUE = 16'h0000)
(
    input clk, resetn,

    // Length of the packets to be output
    output reg[15:0] packet_len,
    
    // How many packets to output
    output reg[31:0] packet_count,
    
    // Number of idle clock-cycles between packets
    output reg[15:0] idle_cycles,

    // Initial value for the first value in the first packet
    output reg[15:0] initial_value,

    // Tells the packet-generator to start generating packets
    output reg start,

    // We use this to reset external logic
    output resetn_out,

    // This is the mismatch alarm that can be raised by the packet checker
    input  alarm,

    // This is asserted when the packet generator is busy generating packets
    input  packet_gen_busy,

    //================== This is an AXI4-Lite slave interface ==================
        
    // "Specify write address"              -- Master --    -- Slave --
    input[AW-1:0]                           S_AXI_AWADDR,   
    input                                   S_AXI_AWVALID,  
    output                                                  S_AXI_AWREADY,
    input[2:0]                              S_AXI_AWPROT,

    // "Write Data"                         -- Master --    -- Slave --
    input[31:0]                             S_AXI_WDATA,      
    input                                   S_AXI_WVALID,
    input[3:0]                              S_AXI_WSTRB,
    output                                                  S_AXI_WREADY,

    // "Send Write Response"                -- Master --    -- Slave --
    output[1:0]                                             S_AXI_BRESP,
    output                                                  S_AXI_BVALID,
    input                                   S_AXI_BREADY,

    // "Specify read address"               -- Master --    -- Slave --
    input[AW-1:0]                           S_AXI_ARADDR,     
    input                                   S_AXI_ARVALID,
    input[2:0]                              S_AXI_ARPROT,     
    output                                                  S_AXI_ARREADY,

    // "Read data back to master"           -- Master --    -- Slave --
    output[31:0]                                            S_AXI_RDATA,
    output                                                  S_AXI_RVALID,
    output[1:0]                                             S_AXI_RRESP,
    input                                   S_AXI_RREADY
    //==========================================================================
);  


//=========================  AXI Register Map  =============================
localparam REG_PACKET_COUNT = 0;
localparam REG_PACKET_LEN   = 1;
localparam REG_IDLE_CYCLES  = 2;
localparam REG_INIT_VALUE   = 3;
localparam REG_BUSY         = 4;
localparam REG_MISMATCH     = 5;
//==========================================================================


//==========================================================================
// Some default values for the registers
//==========================================================================
localparam DEFAULT_PACKET_LEN   = 256;
localparam DEFAULT_IDLE_CYCLES  = 1;
//==========================================================================


//==========================================================================
// We'll communicate with the AXI4-Lite Slave core with these signals.
//==========================================================================
// AXI Slave Handler Interface for write requests
wire[  31:0] ashi_windx;     // Input   Write register-index
wire[AW-1:0] ashi_waddr;     // Input:  Write-address
wire[  31:0] ashi_wdata;     // Input:  Write-data
wire         ashi_write;     // Input:  1 = Handle a write request
reg [   1:0] ashi_wresp;     // Output: Write-response (OKAY, DECERR, SLVERR)
wire         ashi_widle;     // Output: 1 = Write state machine is idle

// AXI Slave Handler Interface for read requests
wire[  31:0] ashi_rindx;     // Input   Read register-index
wire[AW-1:0] ashi_raddr;     // Input:  Read-address
wire         ashi_read;      // Input:  1 = Handle a read request
reg [  31:0] ashi_rdata;     // Output: Read data
reg [   1:0] ashi_rresp;     // Output: Read-response (OKAY, DECERR, SLVERR);
wire         ashi_ridle;     // Output: 1 = Read state machine is idle
//==========================================================================

// The state of the state-machines that handle AXI4-Lite read and AXI4-Lite write
reg ashi_write_state, ashi_read_state;

// The AXI4 slave state machines are idle when in state 0 and their "start" signals are low
assign ashi_widle = (ashi_write == 0) && (ashi_write_state == 0);
assign ashi_ridle = (ashi_read  == 0) && (ashi_read_state  == 0);
   
// These are the valid values for ashi_rresp and ashi_wresp
localparam OKAY   = 0;
localparam SLVERR = 2;
localparam DECERR = 3;

reg[7:0] reset_counter;
assign resetn_out = (resetn == 1) & (reset_counter < 10);

//==========================================================================
// This state machine handles AXI4-Lite write requests
//==========================================================================
always @(posedge clk) begin

    // This strobes high for only a single clock-cycle at a time
    start <= 0;

    // When this is non-zero, resetn_out is asserted
    if (reset_counter) reset_counter <= reset_counter - 1;

    // If we're in reset, initialize important registers
    if (resetn == 0) begin
        reset_counter     <= 0;
        ashi_write_state  <= 0;
        packet_count      <= 0;
        packet_len        <= DEFAULT_PACKET_LEN;
        idle_cycles       <= DEFAULT_IDLE_CYCLES;
        initial_value     <= DEFAULT_INIT_VALUE;

    // Otherwise, we're not in reset...
    end else case (ashi_write_state)
        
        // If an AXI write-request has occured...
        0:  if (ashi_write && !packet_gen_busy) begin
       
                // Assume for the moment that the result will be OKAY
                ashi_wresp <= OKAY;              
            
                // ashi_windex = index of register to be written
                case (ashi_windx)
               
                    REG_PACKET_LEN:
                        if (ashi_wdata > 0 && ashi_wdata <= 9600)
                            packet_len <= ashi_wdata;
                    
                    REG_IDLE_CYCLES:
                        idle_cycles <= ashi_wdata;
                    
                    REG_INIT_VALUE:
                        initial_value <= ashi_wdata;

                    REG_PACKET_COUNT:
                        if (ashi_wdata) begin
                            packet_count     <= ashi_wdata;
                            reset_counter    <= 64;
                            ashi_write_state <= 1;
                         end
                    
 
                    // Writes to any other register are a decode-error
                    default: ashi_wresp <= DECERR;
                endcase
            end

        // Dummy state, doesn't do anything
        1:  if (reset_counter == 0) begin
                start            <= 1;
                ashi_write_state <= 0;
            end

    endcase
end
//==========================================================================





//==========================================================================
// World's simplest state machine for handling AXI4-Lite read requests
//==========================================================================
always @(posedge clk) begin

    // If we're in reset, initialize important registers
    if (resetn == 0) begin
        ashi_read_state <= 0;
    
    // If we're not in reset, and a read-request has occured...        
    end else if (ashi_read) begin
   
        // Assume for the moment that the result will be OKAY
        ashi_rresp <= OKAY;              
        
        // ashi_rindex = index of register to be reads
        case (ashi_rindx)
            
            // Allow a read from any valid register                
            REG_PACKET_LEN:     ashi_rdata <= packet_len;
            REG_PACKET_COUNT:   ashi_rdata <= packet_count;
            REG_IDLE_CYCLES:    ashi_rdata <= idle_cycles;
            REG_INIT_VALUE:     ashi_rdata <= initial_value;
            REG_MISMATCH:       ashi_rdata <= alarm;
            REG_BUSY:           ashi_rdata <= packet_gen_busy;

            // Reads of any other register are a decode-error
            default: ashi_rresp <= DECERR;

        endcase
    end
end
//==========================================================================



//==========================================================================
// This connects us to an AXI4-Lite slave core
//==========================================================================
axi4_lite_slave#(.AW(AW)) i_axi4lite_slave
(
    .clk            (clk),
    .resetn         (resetn),
    
    // AXI AW channel
    .AXI_AWADDR     (S_AXI_AWADDR),
    .AXI_AWPROT     (S_AXI_AWPROT),
    .AXI_AWVALID    (S_AXI_AWVALID),   
    .AXI_AWREADY    (S_AXI_AWREADY),
    
    // AXI W channel
    .AXI_WDATA      (S_AXI_WDATA),
    .AXI_WVALID     (S_AXI_WVALID),
    .AXI_WSTRB      (S_AXI_WSTRB),
    .AXI_WREADY     (S_AXI_WREADY),

    // AXI B channel
    .AXI_BRESP      (S_AXI_BRESP),
    .AXI_BVALID     (S_AXI_BVALID),
    .AXI_BREADY     (S_AXI_BREADY),

    // AXI AR channel
    .AXI_ARADDR     (S_AXI_ARADDR), 
    .AXI_ARPROT     (S_AXI_ARPROT),
    .AXI_ARVALID    (S_AXI_ARVALID),
    .AXI_ARREADY    (S_AXI_ARREADY),

    // AXI R channel
    .AXI_RDATA      (S_AXI_RDATA),
    .AXI_RVALID     (S_AXI_RVALID),
    .AXI_RRESP      (S_AXI_RRESP),
    .AXI_RREADY     (S_AXI_RREADY),

    // ASHI write-request registers
    .ASHI_WADDR     (ashi_waddr),
    .ASHI_WINDX     (ashi_windx),
    .ASHI_WDATA     (ashi_wdata),
    .ASHI_WRITE     (ashi_write),
    .ASHI_WRESP     (ashi_wresp),
    .ASHI_WIDLE     (ashi_widle),

    // ASHI read registers
    .ASHI_RADDR     (ashi_raddr),
    .ASHI_RINDX     (ashi_rindx),
    .ASHI_RDATA     (ashi_rdata),
    .ASHI_READ      (ashi_read ),
    .ASHI_RRESP     (ashi_rresp),
    .ASHI_RIDLE     (ashi_ridle)
);
//==========================================================================



endmodule
